module pd(
  input clock,
  input reset
);
endmodule
