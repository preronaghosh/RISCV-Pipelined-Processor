module register_file #()
(
    
);



endmodule
