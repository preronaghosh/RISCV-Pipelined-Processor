module imemory #()
(
    
);



endmodule
